module ws2812(

);


endmodule